`timescale 1ns / 1ps

module midi_uart_tx_tb;
    // Declare testbench signals

    // Instantiate the DUT
    midi_uart_tx uut (
        // Port mappings
    );

    initial begin
        // Add testbench stimulus
        $finish;
    end

endmodule
