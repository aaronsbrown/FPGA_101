`timescale 1ns / 1ps

module midi_note_sender_tb;
    // Declare testbench signals

    // Instantiate the DUT
    midi_note_sender uut (
        // Port mappings
    );

    initial begin
        // Add testbench stimulus
        $finish;
    end

endmodule
