module flip_flops (
    input clk,
    input rst_n
);

// Add logic here

endmodule
