`timescale 1ns / 1ps

module midi_uart_out_tb;
    // Declare testbench signals

    // Instantiate the DUT
    midi_uart_out uut (
        // Port mappings
    );

    initial begin
        // Add testbench stimulus
        $finish;
    end

endmodule
