module mux_demux (
    input clk,
    input rst_n
);

// Add logic here

endmodule
