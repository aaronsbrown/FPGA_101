`timescale 1ns / 1ps

module seq_player_tb;
    // Declare testbench signals

    // Instantiate the DUT
    seq_player uut (
        // Port mappings
    );

    initial begin
        // Add testbench stimulus
        $finish;
    end

endmodule
