module bpm_clock (
    // Define your module interface here
);
    // Your module implementation goes here
endmodule
