module sequential_logic (
    input clk,
    input rst_n
);

// Add logic here

endmodule
