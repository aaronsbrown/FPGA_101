`timescale 1ns / 1ps

module button_conditioner_tb;
    // Declare testbench signals

    // Instantiate the DUT
    button_conditioner uut (
        // Port mappings
    );

    initial begin
        // Add testbench stimulus
        $finish;
    end

endmodule
