module seq_player (
    // Define your module interface here
);
    // Your module implementation goes here
endmodule
