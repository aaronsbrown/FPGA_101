`timescale 1ns / 1ps

module bpm_clock_tb;
    // Declare testbench signals

    // Instantiate the DUT
    bpm_clock uut (
        // Port mappings
    );

    initial begin
        // Add testbench stimulus
        $finish;
    end

endmodule
