module midi_uart_out (
    // Define your module interface here
);
    // Your module implementation goes here
endmodule
